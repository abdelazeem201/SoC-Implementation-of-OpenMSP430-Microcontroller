
module omsp_multiplier_DW_mult_tc_J3_0 ( a, b, product );
  input [16:0] a;
  input [8:0] b;
  output [25:0] product;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394;
  assign product[25] = 1'b0;
  assign product[24] = 1'b0;

  NBUFFX32 U1 ( .INP(n394), .Z(n1) );
  NBUFFX32 U2 ( .INP(n394), .Z(n2) );
  NBUFFX32 U3 ( .INP(n391), .Z(n3) );
  NBUFFX32 U4 ( .INP(n391), .Z(n4) );
  NBUFFX32 U5 ( .INP(b[2]), .Z(n5) );
  NBUFFX32 U7 ( .INP(n388), .Z(n7) );
  NBUFFX32 U8 ( .INP(n388), .Z(n8) );
  NBUFFX32 U9 ( .INP(n385), .Z(n9) );
  NBUFFX32 U10 ( .INP(n385), .Z(n10) );
  NBUFFX32 U11 ( .INP(n393), .Z(n11) );
  NBUFFX32 U12 ( .INP(n393), .Z(n12) );
  NBUFFX32 U13 ( .INP(n390), .Z(n13) );
  NBUFFX32 U14 ( .INP(n390), .Z(n14) );
  NBUFFX32 U15 ( .INP(b[5]), .Z(n15) );
  NBUFFX32 U17 ( .INP(n387), .Z(n17) );
  NBUFFX32 U18 ( .INP(n387), .Z(n18) );
  NBUFFX32 U19 ( .INP(n384), .Z(n19) );
  NBUFFX32 U20 ( .INP(n384), .Z(n20) );
  NBUFFX32 U21 ( .INP(n392), .Z(n21) );
  NBUFFX32 U22 ( .INP(n392), .Z(n22) );
  NBUFFX32 U23 ( .INP(n389), .Z(n23) );
  NBUFFX32 U24 ( .INP(n389), .Z(n24) );
  NBUFFX32 U25 ( .INP(b[8]), .Z(n25) );
  NBUFFX32 U27 ( .INP(n386), .Z(n27) );
  NBUFFX32 U28 ( .INP(n386), .Z(n28) );
  NBUFFX32 U29 ( .INP(n383), .Z(n29) );
  NBUFFX32 U30 ( .INP(n383), .Z(n30) );
  XOR2X1 U31 ( .IN1(n31), .IN2(n32), .Q(product[23]) );
  XOR2X1 U32 ( .IN1(n55), .IN2(n56), .Q(n31) );
  FADDX1 U33 ( .A(n57), .B(n58), .CI(n33), .CO(n32), .S(product[22]) );
  FADDX1 U34 ( .A(n60), .B(n59), .CI(n34), .CO(n33), .S(product[21]) );
  FADDX1 U35 ( .A(n61), .B(n64), .CI(n35), .CO(n34), .S(product[20]) );
  FADDX1 U36 ( .A(n65), .B(n67), .CI(n36), .CO(n35), .S(product[19]) );
  FADDX1 U37 ( .A(n70), .B(n68), .CI(n37), .CO(n36), .S(product[18]) );
  FADDX1 U38 ( .A(n71), .B(n207), .CI(n38), .CO(n37), .S(product[17]) );
  FADDX1 U39 ( .A(n208), .B(n75), .CI(n39), .CO(n38), .S(product[16]) );
  FADDX1 U40 ( .A(n209), .B(n79), .CI(n40), .CO(n39), .S(product[15]) );
  FADDX1 U41 ( .A(n210), .B(n83), .CI(n41), .CO(n40), .S(product[14]) );
  FADDX1 U42 ( .A(n211), .B(n87), .CI(n42), .CO(n41), .S(product[13]) );
  FADDX1 U43 ( .A(n212), .B(n91), .CI(n43), .CO(n42), .S(product[12]) );
  FADDX1 U44 ( .A(n213), .B(n95), .CI(n44), .CO(n43), .S(product[11]) );
  FADDX1 U45 ( .A(n214), .B(n99), .CI(n45), .CO(n44), .S(product[10]) );
  FADDX1 U46 ( .A(n215), .B(n103), .CI(n46), .CO(n45), .S(product[9]) );
  FADDX1 U47 ( .A(n216), .B(n107), .CI(n47), .CO(n46), .S(product[8]) );
  FADDX1 U48 ( .A(n217), .B(n111), .CI(n48), .CO(n47), .S(product[7]) );
  FADDX1 U49 ( .A(n218), .B(n115), .CI(n49), .CO(n48), .S(product[6]) );
  FADDX1 U50 ( .A(n219), .B(n119), .CI(n50), .CO(n49), .S(product[5]) );
  FADDX1 U51 ( .A(n220), .B(n121), .CI(n51), .CO(n50), .S(product[4]) );
  FADDX1 U52 ( .A(n221), .B(n123), .CI(n52), .CO(n51), .S(product[3]) );
  HADDX1 U53 ( .A0(n222), .B0(n53), .C1(n52), .SO(product[2]) );
  HADDX1 U54 ( .A0(n223), .B0(n54), .C1(n53), .SO(product[1]) );
  HADDX1 U55 ( .A0(n5), .B0(n224), .C1(n54), .SO(product[0]) );
  INVX0 U56 ( .INP(n170), .ZN(n55) );
  INVX0 U57 ( .INP(n56), .ZN(n57) );
  FADDX1 U58 ( .A(n62), .B(n187), .CI(n171), .CO(n58), .S(n59) );
  FADDX1 U59 ( .A(n172), .B(n63), .CI(n188), .CO(n60), .S(n61) );
  INVX0 U60 ( .INP(n62), .ZN(n63) );
  FADDX1 U61 ( .A(n173), .B(n66), .CI(n189), .CO(n64), .S(n65) );
  INVX0 U62 ( .INP(n62), .ZN(n66) );
  FADDX1 U63 ( .A(n69), .B(n72), .CI(n190), .CO(n67), .S(n68) );
  XNOR2X1 U64 ( .IN1(n174), .IN2(n206), .Q(n69) );
  OR2X1 U65 ( .IN1(n174), .IN2(n206), .Q(n62) );
  FADDX1 U66 ( .A(n191), .B(n73), .CI(n74), .CO(n70), .S(n71) );
  HADDX1 U67 ( .A0(n175), .B0(n76), .C1(n72), .SO(n73) );
  FADDX1 U68 ( .A(n192), .B(n77), .CI(n78), .CO(n74), .S(n75) );
  HADDX1 U69 ( .A0(n176), .B0(n80), .C1(n76), .SO(n77) );
  FADDX1 U70 ( .A(n193), .B(n81), .CI(n82), .CO(n78), .S(n79) );
  HADDX1 U71 ( .A0(n177), .B0(n84), .C1(n80), .SO(n81) );
  FADDX1 U72 ( .A(n194), .B(n85), .CI(n86), .CO(n82), .S(n83) );
  HADDX1 U73 ( .A0(n178), .B0(n88), .C1(n84), .SO(n85) );
  FADDX1 U74 ( .A(n195), .B(n89), .CI(n90), .CO(n86), .S(n87) );
  HADDX1 U75 ( .A0(n179), .B0(n92), .C1(n88), .SO(n89) );
  FADDX1 U76 ( .A(n196), .B(n93), .CI(n94), .CO(n90), .S(n91) );
  HADDX1 U77 ( .A0(n180), .B0(n96), .C1(n92), .SO(n93) );
  FADDX1 U78 ( .A(n197), .B(n97), .CI(n98), .CO(n94), .S(n95) );
  HADDX1 U79 ( .A0(n181), .B0(n100), .C1(n96), .SO(n97) );
  FADDX1 U80 ( .A(n198), .B(n101), .CI(n102), .CO(n98), .S(n99) );
  HADDX1 U81 ( .A0(n182), .B0(n104), .C1(n100), .SO(n101) );
  FADDX1 U82 ( .A(n199), .B(n105), .CI(n106), .CO(n102), .S(n103) );
  HADDX1 U83 ( .A0(n183), .B0(n108), .C1(n104), .SO(n105) );
  FADDX1 U84 ( .A(n200), .B(n109), .CI(n110), .CO(n106), .S(n107) );
  HADDX1 U85 ( .A0(n184), .B0(n112), .C1(n108), .SO(n109) );
  FADDX1 U86 ( .A(n201), .B(n113), .CI(n114), .CO(n110), .S(n111) );
  HADDX1 U87 ( .A0(n185), .B0(n116), .C1(n112), .SO(n113) );
  FADDX1 U88 ( .A(n202), .B(n117), .CI(n118), .CO(n114), .S(n115) );
  HADDX1 U89 ( .A0(n25), .B0(n186), .C1(n116), .SO(n117) );
  HADDX1 U90 ( .A0(n203), .B0(n120), .C1(n118), .SO(n119) );
  HADDX1 U91 ( .A0(n204), .B0(n122), .C1(n120), .SO(n121) );
  HADDX1 U92 ( .A0(n15), .B0(n205), .C1(n122), .SO(n123) );
  XOR2X1 U93 ( .IN1(n225), .IN2(n25), .Q(n170) );
  OAI21X1 U94 ( .IN1(n28), .IN2(n337), .IN3(n243), .QN(n225) );
  AOI222X1 U95 ( .IN1(n22), .IN2(n355), .IN3(n24), .IN4(n355), .IN5(n30), 
        .IN6(n358), .QN(n243) );
  XOR2X1 U96 ( .IN1(n226), .IN2(n25), .Q(n56) );
  OAI21X1 U97 ( .IN1(n28), .IN2(n338), .IN3(n244), .QN(n226) );
  AOI222X1 U98 ( .IN1(n22), .IN2(n355), .IN3(n24), .IN4(n358), .IN5(n30), 
        .IN6(n359), .QN(n244) );
  XOR2X1 U99 ( .IN1(n227), .IN2(n25), .Q(n171) );
  OAI21X1 U100 ( .IN1(n28), .IN2(n339), .IN3(n245), .QN(n227) );
  AOI222X1 U101 ( .IN1(n22), .IN2(n358), .IN3(n24), .IN4(n359), .IN5(n30), 
        .IN6(n360), .QN(n245) );
  XOR2X1 U102 ( .IN1(n228), .IN2(n25), .Q(n172) );
  OAI21X1 U103 ( .IN1(n28), .IN2(n340), .IN3(n246), .QN(n228) );
  AOI222X1 U104 ( .IN1(n22), .IN2(n359), .IN3(n24), .IN4(n360), .IN5(n30), 
        .IN6(n361), .QN(n246) );
  XOR2X1 U105 ( .IN1(n229), .IN2(n25), .Q(n173) );
  OAI21X1 U106 ( .IN1(n28), .IN2(n341), .IN3(n247), .QN(n229) );
  AOI222X1 U107 ( .IN1(n22), .IN2(n360), .IN3(n24), .IN4(n361), .IN5(n30), 
        .IN6(n362), .QN(n247) );
  XOR2X1 U108 ( .IN1(n230), .IN2(n25), .Q(n174) );
  OAI21X1 U109 ( .IN1(n28), .IN2(n342), .IN3(n248), .QN(n230) );
  AOI222X1 U110 ( .IN1(n22), .IN2(n361), .IN3(n24), .IN4(n362), .IN5(n30), 
        .IN6(n363), .QN(n248) );
  XOR2X1 U111 ( .IN1(n231), .IN2(n25), .Q(n175) );
  OAI21X1 U112 ( .IN1(n28), .IN2(n343), .IN3(n249), .QN(n231) );
  AOI222X1 U113 ( .IN1(n22), .IN2(n362), .IN3(n24), .IN4(n363), .IN5(n30), 
        .IN6(n364), .QN(n249) );
  XOR2X1 U114 ( .IN1(n232), .IN2(n25), .Q(n176) );
  OAI21X1 U115 ( .IN1(n28), .IN2(n344), .IN3(n250), .QN(n232) );
  AOI222X1 U116 ( .IN1(n22), .IN2(n363), .IN3(n24), .IN4(n364), .IN5(n30), 
        .IN6(n365), .QN(n250) );
  XOR2X1 U117 ( .IN1(n233), .IN2(n25), .Q(n177) );
  OAI21X1 U118 ( .IN1(n28), .IN2(n345), .IN3(n251), .QN(n233) );
  AOI222X1 U119 ( .IN1(n22), .IN2(n364), .IN3(n23), .IN4(n365), .IN5(n29), 
        .IN6(n366), .QN(n251) );
  XOR2X1 U120 ( .IN1(n234), .IN2(n25), .Q(n178) );
  OAI21X1 U121 ( .IN1(n27), .IN2(n346), .IN3(n252), .QN(n234) );
  AOI222X1 U122 ( .IN1(n21), .IN2(n365), .IN3(n23), .IN4(n366), .IN5(n29), 
        .IN6(n367), .QN(n252) );
  XOR2X1 U123 ( .IN1(n235), .IN2(n25), .Q(n179) );
  OAI21X1 U124 ( .IN1(n27), .IN2(n347), .IN3(n253), .QN(n235) );
  AOI222X1 U125 ( .IN1(n21), .IN2(n366), .IN3(n23), .IN4(n367), .IN5(n29), 
        .IN6(n368), .QN(n253) );
  XOR2X1 U126 ( .IN1(n236), .IN2(n25), .Q(n180) );
  OAI21X1 U127 ( .IN1(n27), .IN2(n348), .IN3(n254), .QN(n236) );
  AOI222X1 U128 ( .IN1(n21), .IN2(n367), .IN3(n23), .IN4(n368), .IN5(n29), 
        .IN6(n369), .QN(n254) );
  XOR2X1 U129 ( .IN1(n237), .IN2(n25), .Q(n181) );
  OAI21X1 U130 ( .IN1(n27), .IN2(n349), .IN3(n255), .QN(n237) );
  AOI222X1 U131 ( .IN1(n21), .IN2(n368), .IN3(n23), .IN4(n369), .IN5(n29), 
        .IN6(n370), .QN(n255) );
  XOR2X1 U132 ( .IN1(n238), .IN2(n25), .Q(n182) );
  OAI21X1 U133 ( .IN1(n27), .IN2(n350), .IN3(n256), .QN(n238) );
  AOI222X1 U134 ( .IN1(n21), .IN2(n369), .IN3(n23), .IN4(n370), .IN5(n29), 
        .IN6(n371), .QN(n256) );
  XOR2X1 U135 ( .IN1(n239), .IN2(n25), .Q(n183) );
  OAI21X1 U136 ( .IN1(n27), .IN2(n351), .IN3(n257), .QN(n239) );
  AOI222X1 U137 ( .IN1(n21), .IN2(n370), .IN3(n23), .IN4(n371), .IN5(n29), 
        .IN6(n372), .QN(n257) );
  XOR2X1 U138 ( .IN1(n240), .IN2(n25), .Q(n184) );
  OAI21X1 U139 ( .IN1(n27), .IN2(n352), .IN3(n258), .QN(n240) );
  AOI222X1 U140 ( .IN1(n21), .IN2(n371), .IN3(n23), .IN4(n372), .IN5(n29), 
        .IN6(n373), .QN(n258) );
  XOR2X1 U141 ( .IN1(n241), .IN2(n25), .Q(n185) );
  OAI21X1 U142 ( .IN1(n353), .IN2(n27), .IN3(n259), .QN(n241) );
  INVX0 U143 ( .INP(n124), .ZN(n259) );
  AO22X1 U144 ( .IN1(n21), .IN2(n372), .IN3(n23), .IN4(n373), .Q(n124) );
  XOR2X1 U145 ( .IN1(n242), .IN2(n25), .Q(n186) );
  OAI21X1 U146 ( .IN1(n354), .IN2(n27), .IN3(n260), .QN(n242) );
  INVX0 U147 ( .INP(n125), .ZN(n260) );
  AND2X1 U148 ( .IN1(n21), .IN2(n373), .Q(n125) );
  XNOR2X1 U149 ( .IN1(n261), .IN2(n15), .Q(n187) );
  OAI21X1 U150 ( .IN1(n136), .IN2(n18), .IN3(n280), .QN(n261) );
  AOI222X1 U151 ( .IN1(n12), .IN2(n355), .IN3(n14), .IN4(n355), .IN5(n20), 
        .IN6(n355), .QN(n280) );
  XOR2X1 U152 ( .IN1(n262), .IN2(n15), .Q(n188) );
  OAI21X1 U153 ( .IN1(n18), .IN2(n337), .IN3(n281), .QN(n262) );
  AOI222X1 U154 ( .IN1(n12), .IN2(n355), .IN3(n14), .IN4(n355), .IN5(n20), 
        .IN6(n358), .QN(n281) );
  XOR2X1 U155 ( .IN1(n263), .IN2(n15), .Q(n189) );
  OAI21X1 U156 ( .IN1(n18), .IN2(n338), .IN3(n282), .QN(n263) );
  AOI222X1 U157 ( .IN1(n12), .IN2(n355), .IN3(n14), .IN4(n358), .IN5(n20), 
        .IN6(n359), .QN(n282) );
  XOR2X1 U158 ( .IN1(n264), .IN2(n15), .Q(n190) );
  OAI21X1 U159 ( .IN1(n18), .IN2(n339), .IN3(n283), .QN(n264) );
  AOI222X1 U160 ( .IN1(n12), .IN2(n358), .IN3(n14), .IN4(n359), .IN5(n20), 
        .IN6(n360), .QN(n283) );
  XOR2X1 U161 ( .IN1(n265), .IN2(n15), .Q(n191) );
  OAI21X1 U162 ( .IN1(n18), .IN2(n340), .IN3(n284), .QN(n265) );
  AOI222X1 U163 ( .IN1(n12), .IN2(n359), .IN3(n14), .IN4(n360), .IN5(n20), 
        .IN6(n361), .QN(n284) );
  XOR2X1 U164 ( .IN1(n266), .IN2(n15), .Q(n192) );
  OAI21X1 U165 ( .IN1(n18), .IN2(n341), .IN3(n285), .QN(n266) );
  AOI222X1 U166 ( .IN1(n12), .IN2(n360), .IN3(n14), .IN4(n361), .IN5(n20), 
        .IN6(n362), .QN(n285) );
  XOR2X1 U167 ( .IN1(n267), .IN2(n15), .Q(n193) );
  OAI21X1 U168 ( .IN1(n18), .IN2(n342), .IN3(n286), .QN(n267) );
  AOI222X1 U169 ( .IN1(n12), .IN2(n361), .IN3(n14), .IN4(n362), .IN5(n20), 
        .IN6(n363), .QN(n286) );
  XOR2X1 U170 ( .IN1(n268), .IN2(n15), .Q(n194) );
  OAI21X1 U171 ( .IN1(n18), .IN2(n343), .IN3(n287), .QN(n268) );
  AOI222X1 U172 ( .IN1(n12), .IN2(n362), .IN3(n14), .IN4(n363), .IN5(n20), 
        .IN6(n364), .QN(n287) );
  XOR2X1 U173 ( .IN1(n269), .IN2(n15), .Q(n195) );
  OAI21X1 U174 ( .IN1(n18), .IN2(n344), .IN3(n288), .QN(n269) );
  AOI222X1 U175 ( .IN1(n12), .IN2(n363), .IN3(n14), .IN4(n364), .IN5(n20), 
        .IN6(n365), .QN(n288) );
  XOR2X1 U176 ( .IN1(n270), .IN2(n15), .Q(n196) );
  OAI21X1 U177 ( .IN1(n18), .IN2(n345), .IN3(n289), .QN(n270) );
  AOI222X1 U178 ( .IN1(n12), .IN2(n364), .IN3(n13), .IN4(n365), .IN5(n19), 
        .IN6(n366), .QN(n289) );
  XOR2X1 U179 ( .IN1(n271), .IN2(n15), .Q(n197) );
  OAI21X1 U180 ( .IN1(n17), .IN2(n346), .IN3(n290), .QN(n271) );
  AOI222X1 U181 ( .IN1(n11), .IN2(n365), .IN3(n13), .IN4(n366), .IN5(n19), 
        .IN6(n367), .QN(n290) );
  XOR2X1 U182 ( .IN1(n272), .IN2(n15), .Q(n198) );
  OAI21X1 U183 ( .IN1(n17), .IN2(n347), .IN3(n291), .QN(n272) );
  AOI222X1 U184 ( .IN1(n11), .IN2(n366), .IN3(n13), .IN4(n367), .IN5(n19), 
        .IN6(n368), .QN(n291) );
  XOR2X1 U185 ( .IN1(n273), .IN2(n15), .Q(n199) );
  OAI21X1 U186 ( .IN1(n17), .IN2(n348), .IN3(n292), .QN(n273) );
  AOI222X1 U187 ( .IN1(n11), .IN2(n367), .IN3(n13), .IN4(n368), .IN5(n19), 
        .IN6(n369), .QN(n292) );
  XOR2X1 U188 ( .IN1(n274), .IN2(n15), .Q(n200) );
  OAI21X1 U189 ( .IN1(n17), .IN2(n349), .IN3(n293), .QN(n274) );
  AOI222X1 U190 ( .IN1(n11), .IN2(n368), .IN3(n13), .IN4(n369), .IN5(n19), 
        .IN6(n370), .QN(n293) );
  XOR2X1 U191 ( .IN1(n275), .IN2(n15), .Q(n201) );
  OAI21X1 U192 ( .IN1(n17), .IN2(n350), .IN3(n294), .QN(n275) );
  AOI222X1 U193 ( .IN1(n11), .IN2(n369), .IN3(n13), .IN4(n370), .IN5(n19), 
        .IN6(n371), .QN(n294) );
  XOR2X1 U194 ( .IN1(n276), .IN2(n15), .Q(n202) );
  OAI21X1 U195 ( .IN1(n17), .IN2(n351), .IN3(n295), .QN(n276) );
  AOI222X1 U196 ( .IN1(n11), .IN2(n370), .IN3(n13), .IN4(n371), .IN5(n19), 
        .IN6(n372), .QN(n295) );
  XOR2X1 U197 ( .IN1(n277), .IN2(n15), .Q(n203) );
  OAI21X1 U198 ( .IN1(n17), .IN2(n352), .IN3(n296), .QN(n277) );
  AOI222X1 U199 ( .IN1(n11), .IN2(n371), .IN3(n13), .IN4(n372), .IN5(n19), 
        .IN6(n373), .QN(n296) );
  XOR2X1 U200 ( .IN1(n278), .IN2(n15), .Q(n204) );
  OAI21X1 U201 ( .IN1(n353), .IN2(n17), .IN3(n297), .QN(n278) );
  INVX0 U202 ( .INP(n126), .ZN(n297) );
  AO22X1 U203 ( .IN1(n11), .IN2(n372), .IN3(n13), .IN4(n373), .Q(n126) );
  XOR2X1 U204 ( .IN1(n279), .IN2(n15), .Q(n205) );
  OAI21X1 U205 ( .IN1(n354), .IN2(n17), .IN3(n298), .QN(n279) );
  INVX0 U206 ( .INP(n127), .ZN(n298) );
  AND2X1 U207 ( .IN1(n11), .IN2(n373), .Q(n127) );
  XNOR2X1 U208 ( .IN1(n299), .IN2(n5), .Q(n206) );
  OAI21X1 U209 ( .IN1(n136), .IN2(n8), .IN3(n318), .QN(n299) );
  AOI222X1 U210 ( .IN1(n2), .IN2(n355), .IN3(n4), .IN4(n355), .IN5(n10), .IN6(
        n355), .QN(n318) );
  XOR2X1 U211 ( .IN1(n300), .IN2(n5), .Q(n207) );
  OAI21X1 U212 ( .IN1(n8), .IN2(n337), .IN3(n319), .QN(n300) );
  AOI222X1 U213 ( .IN1(n2), .IN2(n355), .IN3(n4), .IN4(n355), .IN5(n10), .IN6(
        n358), .QN(n319) );
  XOR2X1 U214 ( .IN1(n301), .IN2(n5), .Q(n208) );
  OAI21X1 U215 ( .IN1(n8), .IN2(n338), .IN3(n320), .QN(n301) );
  AOI222X1 U216 ( .IN1(n2), .IN2(n355), .IN3(n4), .IN4(n358), .IN5(n10), .IN6(
        n359), .QN(n320) );
  XOR2X1 U217 ( .IN1(n302), .IN2(n5), .Q(n209) );
  OAI21X1 U218 ( .IN1(n8), .IN2(n339), .IN3(n321), .QN(n302) );
  AOI222X1 U219 ( .IN1(n2), .IN2(n358), .IN3(n4), .IN4(n359), .IN5(n10), .IN6(
        n360), .QN(n321) );
  XOR2X1 U220 ( .IN1(n303), .IN2(n5), .Q(n210) );
  OAI21X1 U221 ( .IN1(n8), .IN2(n340), .IN3(n322), .QN(n303) );
  AOI222X1 U222 ( .IN1(n2), .IN2(n359), .IN3(n4), .IN4(n360), .IN5(n10), .IN6(
        n361), .QN(n322) );
  XOR2X1 U223 ( .IN1(n304), .IN2(n5), .Q(n211) );
  OAI21X1 U224 ( .IN1(n8), .IN2(n341), .IN3(n323), .QN(n304) );
  AOI222X1 U225 ( .IN1(n2), .IN2(n360), .IN3(n4), .IN4(n361), .IN5(n10), .IN6(
        n362), .QN(n323) );
  XOR2X1 U226 ( .IN1(n305), .IN2(n5), .Q(n212) );
  OAI21X1 U227 ( .IN1(n8), .IN2(n342), .IN3(n324), .QN(n305) );
  AOI222X1 U228 ( .IN1(n2), .IN2(n361), .IN3(n4), .IN4(n362), .IN5(n10), .IN6(
        n363), .QN(n324) );
  XOR2X1 U229 ( .IN1(n306), .IN2(n5), .Q(n213) );
  OAI21X1 U230 ( .IN1(n8), .IN2(n343), .IN3(n325), .QN(n306) );
  AOI222X1 U231 ( .IN1(n2), .IN2(n362), .IN3(n4), .IN4(n363), .IN5(n10), .IN6(
        n364), .QN(n325) );
  XOR2X1 U232 ( .IN1(n307), .IN2(n5), .Q(n214) );
  OAI21X1 U233 ( .IN1(n8), .IN2(n344), .IN3(n326), .QN(n307) );
  AOI222X1 U234 ( .IN1(n2), .IN2(n363), .IN3(n4), .IN4(n364), .IN5(n10), .IN6(
        n365), .QN(n326) );
  XOR2X1 U235 ( .IN1(n308), .IN2(n5), .Q(n215) );
  OAI21X1 U236 ( .IN1(n8), .IN2(n345), .IN3(n327), .QN(n308) );
  AOI222X1 U237 ( .IN1(n2), .IN2(n364), .IN3(n3), .IN4(n365), .IN5(n9), .IN6(
        n366), .QN(n327) );
  XOR2X1 U238 ( .IN1(n309), .IN2(n5), .Q(n216) );
  OAI21X1 U239 ( .IN1(n7), .IN2(n346), .IN3(n328), .QN(n309) );
  AOI222X1 U240 ( .IN1(n1), .IN2(n365), .IN3(n3), .IN4(n366), .IN5(n9), .IN6(
        n367), .QN(n328) );
  XOR2X1 U241 ( .IN1(n310), .IN2(n5), .Q(n217) );
  OAI21X1 U242 ( .IN1(n7), .IN2(n347), .IN3(n329), .QN(n310) );
  AOI222X1 U243 ( .IN1(n1), .IN2(n366), .IN3(n3), .IN4(n367), .IN5(n9), .IN6(
        n368), .QN(n329) );
  XOR2X1 U244 ( .IN1(n311), .IN2(n5), .Q(n218) );
  OAI21X1 U245 ( .IN1(n7), .IN2(n348), .IN3(n330), .QN(n311) );
  AOI222X1 U246 ( .IN1(n1), .IN2(n367), .IN3(n3), .IN4(n368), .IN5(n9), .IN6(
        n369), .QN(n330) );
  XOR2X1 U247 ( .IN1(n312), .IN2(n5), .Q(n219) );
  OAI21X1 U248 ( .IN1(n7), .IN2(n349), .IN3(n331), .QN(n312) );
  AOI222X1 U249 ( .IN1(n1), .IN2(n368), .IN3(n3), .IN4(n369), .IN5(n9), .IN6(
        n370), .QN(n331) );
  XOR2X1 U250 ( .IN1(n313), .IN2(n5), .Q(n220) );
  OAI21X1 U251 ( .IN1(n7), .IN2(n350), .IN3(n332), .QN(n313) );
  AOI222X1 U252 ( .IN1(n1), .IN2(n369), .IN3(n3), .IN4(n370), .IN5(n9), .IN6(
        n371), .QN(n332) );
  XOR2X1 U253 ( .IN1(n314), .IN2(n5), .Q(n221) );
  OAI21X1 U254 ( .IN1(n7), .IN2(n351), .IN3(n333), .QN(n314) );
  AOI222X1 U255 ( .IN1(n1), .IN2(n370), .IN3(n3), .IN4(n371), .IN5(n9), .IN6(
        n372), .QN(n333) );
  XOR2X1 U256 ( .IN1(n315), .IN2(n5), .Q(n222) );
  OAI21X1 U257 ( .IN1(n7), .IN2(n352), .IN3(n334), .QN(n315) );
  AOI222X1 U258 ( .IN1(n1), .IN2(n371), .IN3(n3), .IN4(n372), .IN5(n9), .IN6(
        n373), .QN(n334) );
  XOR2X1 U259 ( .IN1(n316), .IN2(n5), .Q(n223) );
  OAI21X1 U260 ( .IN1(n353), .IN2(n7), .IN3(n335), .QN(n316) );
  INVX0 U261 ( .INP(n128), .ZN(n335) );
  AO22X1 U262 ( .IN1(n1), .IN2(n372), .IN3(n3), .IN4(n373), .Q(n128) );
  XOR2X1 U263 ( .IN1(n317), .IN2(n5), .Q(n224) );
  OAI21X1 U264 ( .IN1(n354), .IN2(n7), .IN3(n336), .QN(n317) );
  INVX0 U265 ( .INP(n129), .ZN(n336) );
  AND2X1 U266 ( .IN1(n1), .IN2(n373), .Q(n129) );
  INVX8 U267 ( .INP(n152), .ZN(n337) );
  INVX8 U268 ( .INP(n153), .ZN(n338) );
  INVX8 U269 ( .INP(n154), .ZN(n339) );
  INVX8 U270 ( .INP(n155), .ZN(n340) );
  INVX8 U271 ( .INP(n156), .ZN(n341) );
  INVX8 U272 ( .INP(n157), .ZN(n342) );
  INVX8 U273 ( .INP(n158), .ZN(n343) );
  INVX8 U274 ( .INP(n159), .ZN(n344) );
  INVX8 U275 ( .INP(n160), .ZN(n345) );
  INVX8 U276 ( .INP(n161), .ZN(n346) );
  INVX8 U277 ( .INP(n162), .ZN(n347) );
  INVX8 U278 ( .INP(n163), .ZN(n348) );
  INVX8 U279 ( .INP(n164), .ZN(n349) );
  INVX8 U280 ( .INP(n165), .ZN(n350) );
  INVX8 U281 ( .INP(n166), .ZN(n351) );
  INVX8 U282 ( .INP(n167), .ZN(n352) );
  INVX8 U283 ( .INP(n168), .ZN(n353) );
  INVX8 U284 ( .INP(a[0]), .ZN(n354) );
  NBUFFX4 U285 ( .INP(a[16]), .Z(n355) );
  NBUFFX4 U288 ( .INP(a[15]), .Z(n358) );
  NBUFFX4 U289 ( .INP(a[14]), .Z(n359) );
  NBUFFX4 U290 ( .INP(a[13]), .Z(n360) );
  NBUFFX4 U291 ( .INP(a[12]), .Z(n361) );
  NBUFFX4 U292 ( .INP(a[11]), .Z(n362) );
  NBUFFX4 U293 ( .INP(a[10]), .Z(n363) );
  NBUFFX4 U294 ( .INP(a[9]), .Z(n364) );
  NBUFFX4 U295 ( .INP(a[8]), .Z(n365) );
  NBUFFX4 U296 ( .INP(a[7]), .Z(n366) );
  NBUFFX4 U297 ( .INP(a[6]), .Z(n367) );
  NBUFFX4 U298 ( .INP(a[5]), .Z(n368) );
  NBUFFX4 U299 ( .INP(a[4]), .Z(n369) );
  NBUFFX4 U300 ( .INP(a[3]), .Z(n370) );
  NBUFFX4 U301 ( .INP(a[2]), .Z(n371) );
  NBUFFX4 U302 ( .INP(a[1]), .Z(n372) );
  NBUFFX4 U303 ( .INP(a[0]), .Z(n373) );
  AND3X1 U304 ( .IN1(n374), .IN2(n377), .IN3(n380), .Q(n383) );
  OR2X1 U305 ( .IN1(n374), .IN2(n130), .Q(n386) );
  INVX0 U306 ( .INP(n380), .ZN(n130) );
  AND2X1 U307 ( .IN1(n374), .IN2(n131), .Q(n389) );
  INVX0 U308 ( .INP(n377), .ZN(n131) );
  NOR2X0 U309 ( .IN1(n374), .IN2(n380), .QN(n392) );
  XNOR2X1 U310 ( .IN1(b[6]), .IN2(b[7]), .Q(n377) );
  XNOR2X1 U311 ( .IN1(b[5]), .IN2(b[6]), .Q(n374) );
  XOR2X1 U312 ( .IN1(b[7]), .IN2(b[8]), .Q(n380) );
  AND3X1 U313 ( .IN1(n375), .IN2(n378), .IN3(n381), .Q(n384) );
  OR2X1 U314 ( .IN1(n375), .IN2(n132), .Q(n387) );
  INVX0 U315 ( .INP(n381), .ZN(n132) );
  AND2X1 U316 ( .IN1(n375), .IN2(n133), .Q(n390) );
  INVX0 U317 ( .INP(n378), .ZN(n133) );
  NOR2X0 U318 ( .IN1(n375), .IN2(n381), .QN(n393) );
  XNOR2X1 U319 ( .IN1(b[3]), .IN2(b[4]), .Q(n378) );
  XNOR2X1 U320 ( .IN1(b[2]), .IN2(b[3]), .Q(n375) );
  XOR2X1 U321 ( .IN1(b[4]), .IN2(b[5]), .Q(n381) );
  AND3X1 U322 ( .IN1(n379), .IN2(n382), .IN3(n376), .Q(n385) );
  OR2X1 U323 ( .IN1(n376), .IN2(n134), .Q(n388) );
  INVX0 U324 ( .INP(n382), .ZN(n134) );
  AND2X1 U325 ( .IN1(n376), .IN2(n135), .Q(n391) );
  INVX0 U326 ( .INP(n379), .ZN(n135) );
  NOR2X0 U327 ( .IN1(n382), .IN2(n376), .QN(n394) );
  XNOR2X1 U328 ( .IN1(b[0]), .IN2(b[1]), .Q(n379) );
  INVX0 U329 ( .INP(b[0]), .ZN(n376) );
  XOR2X1 U330 ( .IN1(b[1]), .IN2(b[2]), .Q(n382) );
  INVX0 U331 ( .INP(a[16]), .ZN(n136) );
  FADDX1 U332 ( .A(a[15]), .B(a[16]), .CI(n137), .CO(n152), .S(n153) );
  FADDX1 U333 ( .A(a[14]), .B(a[15]), .CI(n138), .CO(n137), .S(n154) );
  FADDX1 U334 ( .A(a[13]), .B(a[14]), .CI(n139), .CO(n138), .S(n155) );
  FADDX1 U335 ( .A(a[12]), .B(a[13]), .CI(n140), .CO(n139), .S(n156) );
  FADDX1 U336 ( .A(a[11]), .B(a[12]), .CI(n141), .CO(n140), .S(n157) );
  FADDX1 U337 ( .A(a[10]), .B(a[11]), .CI(n142), .CO(n141), .S(n158) );
  FADDX1 U338 ( .A(a[9]), .B(a[10]), .CI(n143), .CO(n142), .S(n159) );
  FADDX1 U339 ( .A(a[8]), .B(a[9]), .CI(n144), .CO(n143), .S(n160) );
  FADDX1 U340 ( .A(a[7]), .B(a[8]), .CI(n145), .CO(n144), .S(n161) );
  FADDX1 U341 ( .A(a[6]), .B(a[7]), .CI(n146), .CO(n145), .S(n162) );
  FADDX1 U342 ( .A(a[5]), .B(a[6]), .CI(n147), .CO(n146), .S(n163) );
  FADDX1 U343 ( .A(a[4]), .B(a[5]), .CI(n148), .CO(n147), .S(n164) );
  FADDX1 U344 ( .A(a[3]), .B(a[4]), .CI(n149), .CO(n148), .S(n165) );
  FADDX1 U345 ( .A(a[2]), .B(a[3]), .CI(n150), .CO(n149), .S(n166) );
  FADDX1 U346 ( .A(a[1]), .B(a[2]), .CI(n151), .CO(n150), .S(n167) );
  HADDX1 U347 ( .A0(a[1]), .B0(a[0]), .C1(n151), .SO(n168) );
endmodule

